--the output is 8-bits, so the INPUT must be 3 bits
